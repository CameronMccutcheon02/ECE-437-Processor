/*
  Cameron McCutcheon

  control unit decode block
*/


module conrol_unit(
    


);


endmodule